`define UNIT_DELAY #1
`define USE_POWER_PINS
`define FUNCTIONAL
`include "libs.ref/sky130_fd_sc_hd/verilog/primitives.v"
`include "libs.ref/sky130_fd_sc_hd/verilog/sky130_fd_sc_hd.v"

